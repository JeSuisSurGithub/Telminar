//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 Education
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Mon Jan 26 19:08:50 2026

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b1;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000FFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_08 = 256'h006666FF66FF6666000000000066666600180000181818180000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h000000000030180C003F6667383C663C00466630180C666200187C063C603E18;
defparam prom_inst_0.INIT_RAM_0A = 256'h000018187E1818000000663CFF3C66000030180C0C0C1830000C18303030180C;
defparam prom_inst_0.INIT_RAM_0B = 256'h006030180C0603000018180000000000000000007E0000003018180000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h003C66061C06663C007E60300C06663C007E181818381818003C6666766E663C;
defparam prom_inst_0.INIT_RAM_0D = 256'h00181818180C667E003C66667C60663C003C6606067C607E0006067F661E0E06;
defparam prom_inst_0.INIT_RAM_0E = 256'h30181800001800000000180000180000003C66063E66663C003C66663C66663C;
defparam prom_inst_0.INIT_RAM_0F = 256'h001800180C06663C0070180C060C18700000007E007E0000000E18306030180E;
defparam prom_inst_0.INIT_RAM_10 = 256'h003C66606060663C007C66667C66667C006666667E663C18003C62606E6E663C;
defparam prom_inst_0.INIT_RAM_11 = 256'h003C66666E60663C006060607860607E007E60607860607E00786C6666666C78;
defparam prom_inst_0.INIT_RAM_12 = 256'h00666C7870786C6600386C0C0C0C0C1E003C18181818183C006666667E666666;
defparam prom_inst_0.INIT_RAM_13 = 256'h003C66666666663C006666666E7E7666006363636B7F7763007E606060606060;
defparam prom_inst_0.INIT_RAM_14 = 256'h003C66063C60663C00666C787C66667C000E3C666666663C006060607C66667C;
defparam prom_inst_0.INIT_RAM_15 = 256'h0063777F6B63636300183C6666666666003C666666666666001818181818187E;
defparam prom_inst_0.INIT_RAM_16 = 256'h003C30303030303C007E6030180C067E001818183C6666660066663C183C6666;
defparam prom_inst_0.INIT_RAM_17 = 256'h7E000000000000000000000000663C18003C0C0C0C0C0C3C0003060C18306000;
defparam prom_inst_0.INIT_RAM_18 = 256'h003C6060603C0000007C66667C606000003E663E063C00000000000000001830;
defparam prom_inst_0.INIT_RAM_19 = 256'h7C063E66663E0000001818183E180E00003C607E663C0000003E66663E060600;
defparam prom_inst_0.INIT_RAM_1A = 256'h00666C786C6060003C06060606000600003C181838001800006666667C606000;
defparam prom_inst_0.INIT_RAM_1B = 256'h003C6666663C000000666666667C000000636B7F7F660000003C181818183800;
defparam prom_inst_0.INIT_RAM_1C = 256'h007C063C603E000000606060667C000006063E66663E000060607C66667C0000;
defparam prom_inst_0.INIT_RAM_1D = 256'h00363E7F6B63000000183C6666660000003E666666660000000E1818187E1800;
defparam prom_inst_0.INIT_RAM_1E = 256'h000E18183018180E007E30180C7E00007C063E666666000000663C183C660000;
defparam prom_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFF0000006E3B000000007018180C1818701818181818181818;
defparam prom_inst_0.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_28 = 256'h00FC62307C30120C00183C60603C180018181818000018000000000000000000;
defparam prom_inst_0.INIT_RAM_29 = 256'h007C063E667C603E181818000018181800187E183C66660000663C66663C6600;
defparam prom_inst_0.INIT_RAM_2A = 256'h0012366C361200000000003E663E063C001C224D514D221C0000000000000066;
defparam prom_inst_0.INIT_RAM_2B = 256'h000000000000003C001C2255595D221C0000000000000000000006067E000000;
defparam prom_inst_0.INIT_RAM_2C = 256'h000000380C180C380000003C30180C38007E18187E18180000000000386C6C38;
defparam prom_inst_0.INIT_RAM_2D = 256'h0000001818000000060606063E66663E607E666666660000000000000000180C;
defparam prom_inst_0.INIT_RAM_2E = 256'h00486C366C4800000000003C6666663C0000003C18183818380C380000000000;
defparam prom_inst_0.INIT_RAM_2F = 256'h003C6660301800180267361C6C3633600762311E2C2663200267361C2C266320;
defparam prom_inst_0.INIT_RAM_30 = 256'h00667E663C186E3B00667E663C18663C00667E663C18180C00667E663C181830;
defparam prom_inst_0.INIT_RAM_31 = 256'h30183C666060663C006F6C6C7E6C3C1F00667E663C3C663C0066667E663C1866;
defparam prom_inst_0.INIT_RAM_32 = 256'h007E6078607E0066007E6078607E663C007E6078607E180C007E6078607E1830;
defparam prom_inst_0.INIT_RAM_33 = 256'h003C1818183C0066003C18183C00663C003C18183C00180C003C18183C001830;
defparam prom_inst_0.INIT_RAM_34 = 256'h003C6666663C180C003C6666663C183000666E7E76666E3B00786C66F6666C78;
defparam prom_inst_0.INIT_RAM_35 = 256'h00663C183C660000003C666666663C66003C6666663C6E3B003C6666663C663C;
defparam prom_inst_0.INIT_RAM_36 = 256'h003C66666600663C003C66666666180C003C666666661830007C66767E6E663E;
defparam prom_inst_0.INIT_RAM_37 = 256'h006C66666C66663C00607C6666667C600018183C6666180C003C666666660066;
defparam prom_inst_0.INIT_RAM_38 = 256'h003E663E063C6E3B003E663E063C663C003E663E063C180C003E663E063C1830;
defparam prom_inst_0.INIT_RAM_39 = 256'h30183C60603C000000376C3F0D3E0000003E66663E3C663C003E663E063C0066;
defparam prom_inst_0.INIT_RAM_3A = 256'h003C607E663C0066003C607E663C663C003C607E663C180C003C607E663C1830;
defparam prom_inst_0.INIT_RAM_3B = 256'h003C181838006600003C18183800663C003C18183800180C003C181838001830;
defparam prom_inst_0.INIT_RAM_3C = 256'h003C6666663C180C003C6666663C183000666666667C6E3B003C66663E060F3C;
defparam prom_inst_0.INIT_RAM_3D = 256'h000018007E001800003C6666663C0066003C6666663C6E3B003C6666663C663C;
defparam prom_inst_0.INIT_RAM_3E = 256'h003E66666666663C003E66666666180C003E666666661830603C6666663C0600;
defparam prom_inst_0.INIT_RAM_3F = 256'h7C063E666666006660607C66667C60007C063E666666180C003E666666660066;

endmodule //Gowin_pROM
