--Copyright (C)2014-2025 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.11.03 Education
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Mon Jan 26 21:22:25 2026

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(10 downto 0)
    );
end Gowin_pROM;

architecture Behavioral of Gowin_pROM is

    signal prom_inst_0_dout_w: std_logic_vector(23 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    dout(7 downto 0) <= prom_inst_0_DO_o(7 downto 0) ;
    prom_inst_0_dout_w(23 downto 0) <= prom_inst_0_DO_o(31 downto 8) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '1',
            BIT_WIDTH => 8,
            RESET_MODE => "ASYNC",
            INIT_RAM_00 => X"00081C3E7F7F7F367EFFE7C3FFDBFF7E7E8199BD81A5817E0000000000000000",
            INIT_RAM_01 => X"0000183C3C1800003E1C3E7F3E1C08083E1C3E7F7F1C3E1C00081C3E7F3E1C08",
            INIT_RAM_02 => X"1E333333BEF0E0F00000000000000000003C664242663C00FFFFE7C3C3E7FFFF",
            INIT_RAM_03 => X"995A3CE7E73C5A990367E6C6C6FEC6FE070F0E0C0CFCCCFC187E183C6666663C",
            INIT_RAM_04 => X"0066006666666666183C7E18187E3C180040707C7F7C70400001071F7F1F0701",
            INIT_RAM_05 => X"FF183C7E187E3C18007E7E7E000000001E331C36361CC67C00D8D8D8DEDBDBFE",
            INIT_RAM_06 => X"00000C067F060C00000018307F30180000183C7E1818181800181818187E3C18",
            INIT_RAM_07 => X"0000183C7EFFFF000000FFFF7E3C180000002466FF66240000007F0303030000",
            INIT_RAM_08 => X"0036367F367F36360000000000363636000C000C0C1E1E0C0000000000000000",
            INIT_RAM_09 => X"0000000000030606006E333B6E1C361C0063660C18336300000C1F301E033E0C",
            INIT_RAM_0A => X"00000C0C3F0C0C000000663CFF3C660000060C1818180C0600180C0606060C18",
            INIT_RAM_0B => X"000103060C183060000C0C0000000000000000003F000000060C0C0000000000",
            INIT_RAM_0C => X"001E33301C30331E003F33061C30331E003F0C0C0C0C0E0C003E676F7B73633E",
            INIT_RAM_0D => X"000C0C0C1830333F001E33331F03061C001E3330301F033F0078307F33363C38",
            INIT_RAM_0E => X"00060C0C000C0C00000C0C00000C0C00000E18303E33331E001E33331E33331E",
            INIT_RAM_0F => X"000C000C1830331E00060C1830180C0600003F00003F000000180C0603060C18",
            INIT_RAM_10 => X"003C66030303663C003F66663E66663F0033333F33331E0C001E037B7B7B633E",
            INIT_RAM_11 => X"007C66730303663C000F06161E16467F007F46161E16467F001F36666666361F",
            INIT_RAM_12 => X"006766361E366667001E333330303078001E0C0C0C0C0C1E003333333F333333",
            INIT_RAM_13 => X"001C36636363361C006363737B6F67630063636B7F7F7763007F66460606060F",
            INIT_RAM_14 => X"001E33380E07331E006766363E66663F00381E3B3333331E000F06063E66663F",
            INIT_RAM_15 => X"0063777F6B636363000C1E3333333333003F333333333333001E0C0C0C0C2D3F",
            INIT_RAM_16 => X"001E06060606061E007F664C1831637F001E0C0C1E3333330063361C1C366363",
            INIT_RAM_17 => X"FF000000000000000000000063361C08001E18181818181E00406030180C0603",
            INIT_RAM_18 => X"001E3303331E0000003B66663E060607006E333E301E00000000000000180C0C",
            INIT_RAM_19 => X"1F303E33336E0000000F06060F06361C001E033F331E0000006E33333E303038",
            INIT_RAM_1A => X"0067361E366606071E33333030300030001E0C0C0C0E000C006766666E360607",
            INIT_RAM_1B => X"001E3333331E000000333333331F000000636B7F7F330000001E0C0C0C0C0C0E",
            INIT_RAM_1C => X"001F301E033E0000000F06666E3B000078303E33336E00000F063E66663B0000",
            INIT_RAM_1D => X"00367F7F6B630000000C1E3333330000006E33333333000000182C0C0C3E0C08",
            INIT_RAM_1E => X"00380C0C070C0C38003F260C193F00001F303E33333300000063361C36630000",
            INIT_RAM_1F => X"007F6363361C08000000000000003B6E00070C0C380C0C070018181800181818",
            INIT_RAM_20 => X"FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3",
            INIT_RAM_21 => X"FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3",
            INIT_RAM_22 => X"FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3",
            INIT_RAM_23 => X"FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3",
            INIT_RAM_24 => X"FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3",
            INIT_RAM_25 => X"FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3",
            INIT_RAM_26 => X"FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3",
            INIT_RAM_27 => X"FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3FFE7FFE7CF9F99C3",
            INIT_RAM_28 => X"003F67060F26361C18187E03037E181800181818180018180000000000000000",
            INIT_RAM_29 => X"1E331C36361CC67C00181818001818180C0C3F0C3F1E333300633E63633E6300",
            INIT_RAM_2A => X"0000CC663366CC0000007E007C36363C7E81B98585B9817E0000000000000063",
            INIT_RAM_2B => X"00000000000000FF7E81A59DA59D817E0000000000000000000030303F000000",
            INIT_RAM_2C => X"0000000E180C180E0000001E060C180E003F000C0C3F0C0C000000001C36361C",
            INIT_RAM_2D => X"000000180000000000D8D8D8DEDBDBFE03063E666666660000000000000C1830",
            INIT_RAM_2E => X"00003366CC66330000003E001C36361C0000001E0C0C0E0C1C30180000000000",
            INIT_RAM_2F => X"001E3303060C000CC3F6ECDF3C66CC07F03366CC7B3363C3C0F3F6ECDB3363C3",
            INIT_RAM_30 => X"00637F63361C3B6E00637F63361C633E0063637F63361C600063637F63361C03",
            INIT_RAM_31 => X"1E30181E3303331E007333337F33367C00333F331E000C0C0063637F63361C63",
            INIT_RAM_32 => X"003F061E063F0033003F061E063F331E003F061E063F0038003F061E063F0007",
            INIT_RAM_33 => X"001E0C0C0C1E0033003C1818183CC37E001E0C0C0C1E0038001E0C0C0C1E0007",
            INIT_RAM_34 => X"001C366363361C60001C366363361C0300333B3F3733003F001F36666F66361F",
            INIT_RAM_35 => X"000063361C36630000183C66663C18C3001C3663361C3B6E001C3663361C633E",
            INIT_RAM_36 => X"003E63636300633E001E333333330038001E333333330007001D36676B73365C",
            INIT_RAM_37 => X"003363331B33331E000F063E663E060F001E0C1E33330038001E333333330033",
            INIT_RAM_38 => X"007E333E301E3B6E00FC667C603CC37E007E333E301E0038007E333E301E0007",
            INIT_RAM_39 => X"1C301E03031E000000FE33FE30FE0000007E333E301E0C0C007E333E301E0033",
            INIT_RAM_3A => X"001E033F331E0033003C067E663CC37E001E033F331E0038001E033F331E0007",
            INIT_RAM_3B => X"001E0C0C0C0E0033003C1818181C633E001E0C0C0C0E001C001E0C0C0C0E0007",
            INIT_RAM_3C => X"001E33331E003800001E33331E000700003333331F001F00001E33333E307E0C",
            INIT_RAM_3D => X"000C0C003F000C0C001E33331E003300001E33331E003B6E001E33331E00331E",
            INIT_RAM_3E => X"007E33333300331E007E333333003800007E333333000700013E676B733E4000",
            INIT_RAM_3F => X"1F303E33330033000F063E66663E06071E303E3333003800007E333333003300"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

end Behavioral; --Gowin_pROM
