--Copyright (C)2014-2025 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.11.03 Education
--Part Number: GW2AR-LV18QN88C8/I7
--Device: GW2AR-18
--Device Version: C
--Created Time: Mon Jan 26 19:52:01 2026

library IEEE;
use IEEE.std_logic_1164.all;

entity Gowin_pROM is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(10 downto 0)
    );
end Gowin_pROM;

architecture Behavioral of Gowin_pROM is

    signal prom_inst_0_dout_w: std_logic_vector(23 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= ad(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    dout(7 downto 0) <= prom_inst_0_DO_o(7 downto 0) ;
    prom_inst_0_dout_w(23 downto 0) <= prom_inst_0_DO_o(31 downto 8) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE => '1',
            BIT_WIDTH => 8,
            RESET_MODE => "SYNC",
            INIT_RAM_00 => X"0010387CFEFEFE6C7EFFE7C3FFDBFF7E7E8199BD81A5817E0000000000000000",
            INIT_RAM_01 => X"0000183C3C1800007C387CFE7C3810107C387CFEFE387C380010387CFE7C3810",
            INIT_RAM_02 => X"78CCCCCC7D0F070F0000000000000000003C664242663C00FFFFE7C3C3E7FFFF",
            INIT_RAM_03 => X"995A3CE7E73C5A99C0E66763637F637FE0F07030303F333F187E183C6666663C",
            INIT_RAM_04 => X"0066006666666666183C7E18187E3C1800020E3EFE3E0E020080E0F8FEF8E080",
            INIT_RAM_05 => X"FF183C7E187E3C18007E7E7E0000000078CC386C6C38633E001B1B1B7BDBDB7F",
            INIT_RAM_06 => X"00003060FE6030000000180CFE0C180000183C7E1818181800181818187E3C18",
            INIT_RAM_07 => X"0000183C7EFFFF000000FFFF7E3C180000002466FF6624000000FEC0C0C00000",
            INIT_RAM_08 => X"006C6CFE6CFE6C6C00000000006C6C6C00300030307878300000000000000000",
            INIT_RAM_09 => X"0000000000C060600076CCDC76386C3800C6663018CCC6000030F80C78C07C30",
            INIT_RAM_0A => X"00003030FC3030000000663CFF3C660000603018181830600018306060603018",
            INIT_RAM_0B => X"0080C06030180C06003030000000000000000000FC0000006030300000000000",
            INIT_RAM_0C => X"0078CC0C380CCC7800FCCC60380CCC7800FC303030307030007CE6F6DECEC67C",
            INIT_RAM_0D => X"00303030180CCCFC0078CCCCF8C060380078CC0C0CF8C0FC001E0CFECC6C3C1C",
            INIT_RAM_0E => X"006030300030300000303000003030000070180C7CCCCC780078CCCC78CCCC78",
            INIT_RAM_0F => X"00300030180CCC78006030180C1830600000FC0000FC000000183060C0603018",
            INIT_RAM_10 => X"003C66C0C0C0663C00FC66667C6666FC00CCCCFCCCCC78300078C0DEDEDEC67C",
            INIT_RAM_11 => X"003E66CEC0C0663C00F06068786862FE00FE6268786862FE00F86C6666666CF8",
            INIT_RAM_12 => X"00E6666C786C66E60078CCCC0C0C0C1E007830303030307800CCCCCCFCCCCCCC",
            INIT_RAM_13 => X"00386CC6C6C66C3800C6C6CEDEF6E6C600C6C6D6FEFEEEC600FE6662606060F0",
            INIT_RAM_14 => X"0078CC1C70E0CC7800E6666C7C6666FC001C78DCCCCCCC7800F060607C6666FC",
            INIT_RAM_15 => X"00C6EEFED6C6C6C6003078CCCCCCCCCC00FCCCCCCCCCCCCC007830303030B4FC",
            INIT_RAM_16 => X"007860606060607800FE6632188CC6FE0078303078CCCCCC00C66C38386CC6C6",
            INIT_RAM_17 => X"FF0000000000000000000000C66C381000781818181818780002060C183060C0",
            INIT_RAM_18 => X"0078CCC0CC78000000DC66667C6060E00076CC7C0C7800000000000000183030",
            INIT_RAM_19 => X"F80C7CCCCC76000000F06060F0606C380078C0FCCC7800000076CCCC7C0C0C1C",
            INIT_RAM_1A => X"00E66C786C6660E078CCCC0C0C0C000C007830303070003000E66666766C60E0",
            INIT_RAM_1B => X"0078CCCCCC78000000CCCCCCCCF8000000C6D6FEFECC00000078303030303070",
            INIT_RAM_1C => X"00F80C78C07C000000F0606676DC00001E0C7CCCCC760000F0607C6666DC0000",
            INIT_RAM_1D => X"006CFEFED6C60000003078CCCCCC00000076CCCCCCCC000000183430307C3010",
            INIT_RAM_1E => X"001C3030E030301C00FC643098FC0000F80C7CCCCCCC000000C66C386CC60000",
            INIT_RAM_1F => X"00FEC6C66C381000000000000000DC7600E030301C3030E00018181800181818",
            INIT_RAM_20 => X"FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3",
            INIT_RAM_21 => X"FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3",
            INIT_RAM_22 => X"FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3",
            INIT_RAM_23 => X"FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3",
            INIT_RAM_24 => X"FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3",
            INIT_RAM_25 => X"FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3",
            INIT_RAM_26 => X"FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3",
            INIT_RAM_27 => X"FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3FFE7FFE7F3F999C3",
            INIT_RAM_28 => X"00FCE660F0646C3818187EC0C07E181800181818180018180000000000000000",
            INIT_RAM_29 => X"78CC386C6C38633E00181818001818183030FC30FC78CCCC00C67CC6C67CC600",
            INIT_RAM_2A => X"00003366CC66330000007E003E6C6C3C7E819DA1A19D817E00000000000000C6",
            INIT_RAM_2B => X"00000000000000FF7E81A5B9A5B9817E000000000000000000000C0CFC000000",
            INIT_RAM_2C => X"0000007018301870000000786030187000FC003030FC303000000000386C6C38",
            INIT_RAM_2D => X"0000001800000000001B1B1B7BDBDB7FC0607C6666666600000000000030180C",
            INIT_RAM_2E => X"0000CC663366CC0000007C00386C6C380000007830307030380C180000000000",
            INIT_RAM_2F => X"0078CCC060300030C36F37FB3C6633E00FCC6633DECCC6C303CF6F37DBCCC6C3",
            INIT_RAM_30 => X"00C6FEC66C38DC7600C6FEC66C38C67C00C6C6FEC66C380600C6C6FEC66C38C0",
            INIT_RAM_31 => X"780C1878CCC0CC7800CECCCCFECC6C3E00CCFCCC7800303000C6C6FEC66C38C6",
            INIT_RAM_32 => X"00FC607860FC00CC00FC607860FCCC7800FC607860FC001C00FC607860FC00E0",
            INIT_RAM_33 => X"00783030307800CC003C1818183CC37E007830303078001C00783030307800E0",
            INIT_RAM_34 => X"00386CC6C66C380600386CC6C66C38C000CCDCFCECCC00FC00F86C66F6666CF8",
            INIT_RAM_35 => X"0000C66C386CC60000183C66663C18C300386CC66C38DC7600386CC66C38C67C",
            INIT_RAM_36 => X"007CC6C6C600C67C0078CCCCCCCC001C0078CCCCCCCC00E000B86CE6D6CE6C3A",
            INIT_RAM_37 => X"00CCC6CCD8CCCC7800F0607C667C60F000783078CCCC001C0078CCCCCCCC00CC",
            INIT_RAM_38 => X"007ECC7C0C78DC76003F663E063CC37E007ECC7C0C78001C007ECC7C0C7800E0",
            INIT_RAM_39 => X"380C78C0C0780000007FCC7F0C7F0000007ECC7C0C783030007ECC7C0C7800CC",
            INIT_RAM_3A => X"0078C0FCCC7800CC003C607E663CC37E0078C0FCCC78001C0078C0FCCC7800E0",
            INIT_RAM_3B => X"00783030307000CC003C18181838C67C007830303070003800783030307000E0",
            INIT_RAM_3C => X"0078CCCC78001C000078CCCC7800E00000CCCCCCF800F8000078CCCC7C0C7E30",
            INIT_RAM_3D => X"00303000FC0030300078CCCC7800CC000078CCCC7800DC760078CCCC7800CC78",
            INIT_RAM_3E => X"007ECCCCCC00CC78007ECCCCCC001C00007ECCCCCC00E000807CE6D6CE7C0200",
            INIT_RAM_3F => X"F80C7CCCCC00CC00F0607C66667C60E0780C7CCCCC001C00007ECCCCCC00CC00"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

end Behavioral; --Gowin_pROM
